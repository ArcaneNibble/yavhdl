type test is access bar foo (baz'range);
