architecture aaa of bbb(ccc).ddd is
    signal foo : bar;
    signal baz : qux;
begin
    asdf <= fdsa;
end architecture eee;
