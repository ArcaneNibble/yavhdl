foo(bar range 0 to 2)