type foo is (a, b, c, d);
