entity test is
    type t is protected body end protected;
end;
