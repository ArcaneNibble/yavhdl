entity test is
    subtype t is baz."=" foo'bar;
end;
