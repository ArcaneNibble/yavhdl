entity test is
    type test is (foo, foo);
begin end;
