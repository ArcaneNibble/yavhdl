entity 0test is end;
