entity test is
    file foo : bar open qux is "baz";
end;
