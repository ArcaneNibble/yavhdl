[foo, bar, baz, qux return asdf]