new STRING (1 to 10)(2 to 11)