architecture test of test2 is
    constant foo : bar := "hello";
begin end;
