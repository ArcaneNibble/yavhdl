entity test is
    constant a : b :=
    foo'(bar, baz|others => qux);
end;
