entity test is
    constant a : b :=
    foo(5).bar;
end;
