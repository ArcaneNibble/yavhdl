process
    type t is protected body
        procedure p;
    end protected body u;
begin
end process;
