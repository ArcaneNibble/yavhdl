use foo.bar;
entity test is end;
