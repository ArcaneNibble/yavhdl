configuration xxx of xxx is
    for xxx
        for aaa : bbb
            generic map (ccc => ddd);
            use vunit a;
            for yyy
            end for;
        end for;
    end for;
end configuration xxx;
