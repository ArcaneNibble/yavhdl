process
    procedure aaa is new bbb generic map(
        zzz => iii(jjj(
            foo1(bar range baz'qux)(open),
            foo2(bar range baz'qux)
        ))
    );
begin
end process;
