5 ns
