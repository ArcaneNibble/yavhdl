entity test is
    type t is range 2 downto 0;
end;
