architecture a of a is begin
   result <= foo(bar => 3, baz => 4)(3);
end;
