library foo;
entity test is end;
