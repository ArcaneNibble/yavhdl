a * b + c