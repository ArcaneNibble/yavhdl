postponed with asdf select a <= b when c, d when e;
