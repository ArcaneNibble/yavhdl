<<constant foo : baz bar>>