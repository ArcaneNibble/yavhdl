entity test is
    constant a : b :=
    foo /= bar nand baz nor qux;
end;
