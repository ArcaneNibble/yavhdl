process
    type t is protected
        procedure p;
    end protected u;
begin
end process;
