'a'.'b''c."e"'f