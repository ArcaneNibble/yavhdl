process
    procedure foo (
        procedure aaa;
        procedure bbb is <>;
        procedure ccc is ddd
    );
begin
end process;
