entity test is
    constant a : b :=
    new foo'(bar);
end;
