l: block
    for a : b;
begin end block;
