if 123 then
    foo(aaa, bbb, ccc, ddd, open, eee, fff => ggg, hhh, iii, open, bar.baz.qux."wat"(jjj) => open, kkk);
end if;
