architecture test of test2 is
    signal foo : bar := baz;
begin end;
