entity test is
    constant a : b :=
    foo(0 to 2)'bar(bax);
end;
