entity test is
    type t is file of foo;
end;
