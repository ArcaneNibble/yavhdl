entity test is
    type t is record
    end record;
end;
