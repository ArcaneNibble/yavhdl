entity test is
    subtype t is foo(bar (open)(open));
end;
