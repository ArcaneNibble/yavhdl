entity test is
    type foo is (foo, bar);
    --type test is ('a', 'b');
    type testtype is (foo, bar);
    type foo is (baz);
begin end;
