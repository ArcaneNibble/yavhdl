mylabel: entity foo(bar).baz(qux);
