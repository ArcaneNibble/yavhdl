entity test is end;
