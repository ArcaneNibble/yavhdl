foo(bar (0 to 2))