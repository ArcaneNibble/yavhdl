entity test is
    package a is new b generic map(foo, open, bar);
end;
