 entity test is begin end;
entity test is begin end;
entity \test3\ is begin end;
