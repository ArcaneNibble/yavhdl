entity test is
    file foo : bar is "baz";
end;
