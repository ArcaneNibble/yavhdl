entity test is
    type t is array(0 to 1, 2 to 3) of foo;
end;
