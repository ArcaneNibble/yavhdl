foo(bar (0 to 2, 1 to 3, 2 to 4, 3 to 5)(baz (111 to 222)))