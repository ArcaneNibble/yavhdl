entity test is
    subtype t is ((bar baz, qux zzz)) foo;
end;
