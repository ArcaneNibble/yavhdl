entity test is
    constant a : b :=
    <<constant foo : t>>;
end;
