entity \test
\ is end;
