entity test is
    subtype t is foo'subtype range bar'baz;
end;
