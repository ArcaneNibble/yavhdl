configuration aaa of bbb is
    use a.b;
    use vunit c;

    for xxx(yyy).zzz(www range iii'jjj)
    end for;
end configuration ccc;
