type foo is range 0 to 5;
