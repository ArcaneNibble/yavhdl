process
    procedure foo generic map(
        aaa => bbb,
        ccc(ddd) => inertial eee
    );
begin
end process;
