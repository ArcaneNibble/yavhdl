architecture test of test2 is
    constant foo : bar;
begin end;
