postponed a <= guarded transport b;
