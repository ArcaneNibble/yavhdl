entity test is
    type t is array(0 to 2, tt range <>) of foo;
end;
