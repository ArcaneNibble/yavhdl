process
    package aaa is new bbb;
    package ccc is new ddd generic map(ggg(eee) => hhh(fff, ggg, bar range baz'qux)(0 to 2, 1 to 3));
begin
end process;
