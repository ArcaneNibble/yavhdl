entity test is
    type test1 is (foo);
    constant test2, test3 : test1;
begin end;
