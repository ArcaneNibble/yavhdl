process
    procedure aaa is new bbb [] generic map (ccc);
begin
end process;
