entity test is
    package a is new b generic map(c => ((bar baz, qux zzz)) foo);
end;
