entity test is
    type t is range 0 to 1e2;
end;
