process
    group aaa : bbb(ddd, eee, fff'ggg'hhh, "iii", "jjj", kkk(lll));
begin
end process;
