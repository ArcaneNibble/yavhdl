process
    procedure p generic(
        package aaa is new bbb generic map(default)
    );
begin
end process;
