entity test is
    type t is record
        foo, bar : baz;
    end record;
end;
