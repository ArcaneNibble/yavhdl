entity test is
    type test is (foo);
    function test1 (constant a : test) return test;
begin end;
