entity test is
    type t;
end;
