process
    procedure foo generic map(
    );
begin
end process;
