entity test is
    type t is range 0 to 1.e2;
end;
