entity test is--This is a comment a��������������������
end;
