entity test is
    type t is array(0 to 1) of foo;
end;
