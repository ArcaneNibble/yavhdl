foo(

bar

(baz (0 to 2), qux (1 to 3))

)