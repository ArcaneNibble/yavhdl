entity test is
    type t is range 0 to 16#g.f#2;
end;
