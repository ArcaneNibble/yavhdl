entity test is
    subtype t is foo(open)(open);
end;
