type test is record
    aaa,bbb,ccc : bar foo (baz'range);
    ddd: eee;
end record;
