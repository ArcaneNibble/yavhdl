with asdf select? (foo, bar, baz, a|b|c|d => qux) <= force out
    aaa when 111,
    bbb when 222;
