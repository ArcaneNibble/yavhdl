\������������������������������\
