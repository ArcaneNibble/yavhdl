architecture test of test2 is
    constant foo : bar := 32X"12345";
begin end;
