entity test is
    type test is (foo);
    type test is (bar);
begin end;
