with asdf select? foo :=
    aaa when 111,
    bbb when 222,
    zzz when others;
