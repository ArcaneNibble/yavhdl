entity test is
    --type foo is (foo, bar);
    type test is ('a', 'a');
    type testtype is (foo, bar);
    --type foo is (baz);
begin end;
