entity test is
    type t is range foo'bar;
end;
