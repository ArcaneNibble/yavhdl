entity test is
    constant a : b :=
    foo(5)(0 to 2);
end;
