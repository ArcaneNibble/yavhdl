context foo.bar;
entity test is end;
