process
    attribute aaa : bbb;
begin
end process;
