process
    attribute aaa of bbb [], ccc, "ddd", 'e' [fff, ggg return hhh]: property is zzz;
begin
end process;
