entity test is
    type t is range 0 to 1E-2;
end;
