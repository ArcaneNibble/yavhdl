process
    file aaa,bbb : ccc;
    file ddd,eee : fff is ggg;
    file hhh,iii : jjj open kkk is lll;

    alias mmm is nnn;
    alias ooo : ppp is qqq;
    alias "rrr" : sss is ttt [uuu, vvv return www];
begin
end process;
