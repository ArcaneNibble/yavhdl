foo((((((((((((bar))))))))))) baz)