entity test is
    subtype t is bar foo'subtype range 0 to 2;
end;
