entity test is
    constant a : b :=
    (a + b) * c;
end;
