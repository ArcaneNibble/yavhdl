architecture test of test2 is
    constant foo, foo2 : bar := baz;
begin end;
