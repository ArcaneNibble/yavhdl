foo(bar baz)