context aaa is
    library a, b;
end;
