entity test is
    subtype t is foo;
end;
