architecture test of test2 is
    constant foo : bar := 32sO"12345";
begin end;
