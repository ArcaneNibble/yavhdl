context foo;
entity test is end;
