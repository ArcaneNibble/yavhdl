(foo, baz) <= reject 123 ps inertial null after 10 ns, 123 after 20 ns;