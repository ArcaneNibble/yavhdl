process
    procedure foo (
        file aaa : bbb;
        ccc : ddd;
        eee : fff := ggg;
        hhh : inout iii;
        jjj : linkage kkk := lll
    );
begin
end process;
