entity test is
    constant a : b :=
    <<constant @foo.bar.baz : t>>;
end;
