architecture test of test2 is begin end;