entity test is
    constant a : b :=
    foo'(bar, aa+bb|cc'dd => qux);
end;
