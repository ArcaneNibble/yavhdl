architecture test of test2 is
    shared variable foo, foo2 : bar := baz;
begin end;
