process
begin
    foo <= bar;
    baz <= qux;
end;
