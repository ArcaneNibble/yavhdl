

foo -- single line comment
bar

/* comment with

multiple

/*

lines */


�
