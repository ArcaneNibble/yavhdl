mylabel: postponed asdf(fdsa, aaa => bbb);
