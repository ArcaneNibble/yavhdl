entity test is/*This is a /*comment*/end;
