with asdf select? (foo, bar, baz, a|b|c|d => qux) <= reject 666 inertial
    aaa, zzz when 111,
    bbb when 222;
