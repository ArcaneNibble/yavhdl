entity test is
    constant a : b :=
    ??foo;
end;
