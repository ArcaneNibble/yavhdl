entity test is begin end;
entity test2 is begin end;
entity \test3\ is begin end;
