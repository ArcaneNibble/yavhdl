foo(aaa, bbb, ccc, ddd, open, eee, fff => ggg, hhh, iii, open, jjj => open, kkk)