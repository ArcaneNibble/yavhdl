<<constant foo : bar>>