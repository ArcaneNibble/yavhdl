architecture test of test2 is
    constant foo : bar := "hel"lo";
begin end;
