process
    attribute aaa of bbb:property is ccc;
begin
end process;
