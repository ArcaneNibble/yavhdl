mylabel: block

generic(aaa : bbb);
generic map(ccc => ddd);
port(xxx : yyy);
port map(zzz => www);

begin end block;
