entity test is
    constant a : b :=
    <<constant foo(bar) : t>>;
end;
