12UB"X1"