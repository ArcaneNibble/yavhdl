package test is
    subtype test2 is test1;
end;
