architecture test of test2 is
    constant foo : bar := 32o"12345";
begin end;
