process
    package p is
        disconnect others:zzz after 5 ns;
    end;
begin
end process;
