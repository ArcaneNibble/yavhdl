foo.all ** bar.baz
