foo(asdf range bar'baz(qux))