process
    procedure foo (
        aaa : bbb bus;
        ccc : inout ddd bus;
        eee : fff bus := ggg;
        hhh : linkage iii bus := jjj
    );
begin
end process;
