foo'bar(baz)