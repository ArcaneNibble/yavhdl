with asdf select? foo :=
    aaa'range when 111,
    bbb'subtype when 222,
    zzz when others;
