entity test begin end;
