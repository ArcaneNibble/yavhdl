entity test is
    function test1 return test;
    impure function test2 return test;
begin end;
