entity test is
    package a is new b generic map(c => foo'subtype range bar'baz);
end;
