mylabel: configuration foo(bar).baz(qux).zzz generic map (aaa) port map (bbb);
