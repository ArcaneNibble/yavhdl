postponed with asdf select? a guarded transport <= b when c, d when e;
postponed with asdf select? a guarded transport <= b when c, d when e;
