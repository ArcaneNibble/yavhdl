entity test is
    subtype t is foo'subtype range 0 to 2;
end;
