entity test is
    type test is (foo);
    function test1 (a : test) return test;
begin end;
