(foo, aaa|bbb|ccc'ddd(eee) => bar)