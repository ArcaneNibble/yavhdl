entity test is
    subtype t is foo'bar;
end;
