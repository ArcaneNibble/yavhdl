entity test is
    constant a : b :=
    new foo;
end;
