configuration aaa of bbb is
    use a.b;
    use vunit c;
end configuration ccc;
