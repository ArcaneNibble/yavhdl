entity test� is end;
