entity test is begin end;
