entity test is
    subtype t is ((bar)) foo;
end;
