package foo is new bar;
