entity test is begin end;
entity test is begin end;
