entity \test\ is end;
