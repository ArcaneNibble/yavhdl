entity \/*this isn't a comment*/\ is end;
