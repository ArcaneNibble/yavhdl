entity test is
    constant a : b :=
    foo /= bar nand nand baz;
end;
