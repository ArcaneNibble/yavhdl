entity test is
    type t is (foo, bar, 'b', 'q');
end;
