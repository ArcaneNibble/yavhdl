entity test is
    subtype t is ((bar baz)) foo;
end;
