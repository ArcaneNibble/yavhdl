architecture test of test2 is
    constant foo : bar := 32d"12345";
begin end;
