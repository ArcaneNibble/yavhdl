foo(open, zzz, qux => asdf, bar => baz'aaa(bbb))