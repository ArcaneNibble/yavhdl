architecture test of test2 is
    signal foo, foo2 : bar := baz;
begin end;
