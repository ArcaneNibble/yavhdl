entity test is
    subtype t is foo range bar'baz;
end;
