if 123 then
    foo(aaa, bbb, ccc, ddd, open, eee, fff => ggg, hhh, iii, open, bar.baz.qux."wat"(jjj) => open, kkk);
elsif 456 then
    bar(111);
elsif 789 then
else
    baz(222);
end if mylabel;
