process
    procedure aaa is
        procedure bbb is begin end function bbb;
    begin
        xxx <= yyy;
    end procedure zzz;
begin
end process;
