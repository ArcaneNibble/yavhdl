architecture test of test2 is
    constant foo : bar := baz;
begin end;
