entity test is
    constant a : b :=
    foo + bar;
end;
