l: case zzz generate
    when a =>
    when b =>
end generate l2;
