architecture test of test2 is
    variable foo : bar := baz;
begin end;
