entity test is
    subtype t is foo(bar)(0 to 2);
end;
