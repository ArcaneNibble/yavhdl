entity test is
    subtype t is foo(open)(bar);
end;
