process
    use x.y;
    use z.all;
    use a.b, c.d, e.f;
begin
end process;
