(foo, bar, baz, qux)