entity test is
    type test is (foo);
    function test1 return test;
    impure function test2 return test;
begin end;
