entity test is
    type t is range 0 to 1.0.E+2;
end;
