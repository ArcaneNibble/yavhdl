process
    group aaa is (signal);
    group bbb is (signal, label);
    group ccc is (signal<>);
    group ccc is (signal<>, label);
    group ccc is (signal<>, label<>);
begin
end process;
