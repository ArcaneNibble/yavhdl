entity test is
    package a is new b generic map(c => baz foo'bar);
end;
