process
    package body test is
        package body aaa is end;
        package body bbb is end package body;
        package body ccc is end ddd;
        package body eee is end package body fff;
    end;
begin
end process;
