package body test is end;
