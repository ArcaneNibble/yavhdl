(foo, bar, baz, a|b|c|d => qux) <= reject 666 inertial
    aaa when 111
    else bbb when 222
    else ccc when 333
    else ddd;
