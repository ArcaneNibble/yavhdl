foo(


base range foo'bar


)