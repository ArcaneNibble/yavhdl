package test is end;
