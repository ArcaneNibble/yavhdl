entity test is
    subtype t is foo(bar (open)(baz (quz'xxx)));
end;
