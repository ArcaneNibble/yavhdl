entity test is
    type t is array(tt range <>) of foo;
end;
