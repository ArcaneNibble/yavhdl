postponed a <= b;
