l: block
    for others : z
        use entity aaa(bbb).ccc(ddd)
        generic map(eee => fff)
        port map(ggg => hhh)
    ;
begin end block;
