l: if aaa: 1 generate
elsif 2 generate
elsif bbb: 3 generate
else zzz: generate
end generate l2;
