process
    procedure foo generic map(
        (x."bbb") ccc (ddd)
    );
begin
end process;
