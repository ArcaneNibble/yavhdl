type asdf is array (aaa range <>, bbb range <>) of bar foo (baz'range);