process
    procedure aaa generic();
    procedure bbb generic() ();
    procedure ccc generic() parameter ();
    function ddd generic() return zzz;
    function eee generic() () return zzz;
    function fff generic() parameter () return zzz;
begin
end process;
