process
    package test is generic(xxx:yyy); generic map (aaa => bbb); 
        package aaa is end;
        package bbb is end package;
        package ccc is end ddd;
        package eee is end package fff;
    end;
begin
end process;
