process
    procedure foo generic map(
        aaa => x."bbb" ccc
    );
begin
end process;
