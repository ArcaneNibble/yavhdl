foo.all
