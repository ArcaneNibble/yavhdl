type test is file of string;
