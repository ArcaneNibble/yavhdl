case? 123 is
    when 1|2 =>
        foo(bar);
    when 4 to 10 =>
        baz(qux);
    when your'mom =>
    when others =>
end case? mylabel;
