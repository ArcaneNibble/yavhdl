entity zzz is
    generic(aaa:bbb);
    port(ccc:ddd);
begin
    assert a;
end;
