entity test is begin end;
entity test2 is begin end test5;
entity \test3\ is begin end;
