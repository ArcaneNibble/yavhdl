entity test is
    constant a : b :=
    null;
end;
