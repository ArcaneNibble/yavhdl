foo(bar(baz (asdf'fdsa(123)), qux (1 to 3)))