label1: postponed process--(xxx, yyy, zzz)
    type aaa is range 0 to 5;
    type bbb is range 5 to 10;
begin
    foo <= bar;
    baz <= qux;
end postponed process label2;
