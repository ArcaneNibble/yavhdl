mylabel: component foo;
