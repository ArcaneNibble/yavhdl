entity test is
    type t is access foo;
end;
