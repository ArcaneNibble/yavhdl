process
    procedure aaa is new bbb generic map(
        zzz => foo(bar, baz)
    );
begin
end process;
