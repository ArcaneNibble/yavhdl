process
    package aaa is new bbb;
    package ccc is new ddd generic map(ggg(eee) => hhh(open)(open));
begin
end process;
