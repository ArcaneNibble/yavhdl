architecture test of test2 is
    constant foo : bar := 32b"12345";
begin end;
