entity test is
    file foo : bar;
end;
