foo(


(a b, c d, e f, g (h i)) base


)