entity test is
    subtype test is test;
begin end;
