mylabel: postponed assert asdf(fdsa, aaa => bbb);
