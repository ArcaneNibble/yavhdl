l: block
    for others : z;
        use vunit a, b, c;
        use vunit d;
    end for;
begin end block;
