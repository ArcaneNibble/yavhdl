entity test is
    type t is file foo;
end;
