16#E#E1