entity _test is end;
