foo(bar, baz, qux)