main_name[foo, bar, baz, qux return asdf]'attrib(arg1 + arg2)