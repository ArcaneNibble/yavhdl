for asdf in 0 to 2 loop
    foo(bar);
    baz(qux);
end loop mylabel;
