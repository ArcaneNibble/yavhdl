entity test is
    subtype t is foo(open);
end;
