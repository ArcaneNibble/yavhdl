process
    package aaa is new bbb;
    package ccc is new ddd generic map(ggg(eee) => hhh(fff, ggg, bar range baz'qux)(open));
begin
end process;
