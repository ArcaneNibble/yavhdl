process
    procedure foo (
        function aaa return xxx;
        pure function bbb return yyy;
        impure function ccc return zzz;

        function ddd (eee : fff) return ggg;
        function hhh parameter (iii : jjj) return kkk
    );
begin
end process;
