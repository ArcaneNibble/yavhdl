(foo, baz) <= release in;