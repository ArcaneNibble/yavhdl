entity test_ is end;
