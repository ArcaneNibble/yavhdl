entity test is
    package a is new b generic map(inertial foo);
end;
