entity test is
    type t is protected end protected;
end;
