architecture test of test2 is
    constant foo : bar := 32Ub"12345";
begin end;
