context test is end;
