use foo;
entity test is end;
