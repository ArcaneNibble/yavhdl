entity test is
    type test1 is (foo, bar);
    type test2 is (foo, baz);
begin end;
