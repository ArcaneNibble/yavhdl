architecture test of foo.bar.baz.qux is begin end;