entity test is begin end;
entity test2 is begin end;
