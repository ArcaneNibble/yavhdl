entity test is
    type t is range 0 to 2#1.1#2;
end;
