entity test is
    subtype t is foo(0 to 2)(bar);
end;
