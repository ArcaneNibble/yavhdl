entity test is
    package a is new b generic map(bar(baz) => inertial foo);
end;
