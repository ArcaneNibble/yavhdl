process
    procedure aaa;
    procedure bbb (file xxx : yyy; file vvv : www);
    procedure ccc parameter (file xxx : yyy);
    function ddd return zzz;
    function eee (file xxx : yyy) return zzz;
    function fff parameter (file xxx : yyy) return zzz;
begin
end process;
