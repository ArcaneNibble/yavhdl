<<constant foo : bar baz (qux (0 to 2), asdf (fdsa (open)(0 to 2)))>>