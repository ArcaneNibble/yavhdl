entity \t\\est\ is end;
