(foo, baz) <= null after 10 ns, 123 after 20 ns;