entity test is
    type test is (foo);
begin end;
