process
    procedure foo;
begin
end process;
