entity test is
    file foo : bar open qux;
end;
