process
    procedure aaa is new bbb generic map(
        zzz => foo(bar (open)(open))
    );
begin
end process;
