process
    procedure aaa is new bbb generic map(
        zzz => iii(jjj(
            foo(bar range baz'qux)(open)
        ))
    );
begin
end process;
