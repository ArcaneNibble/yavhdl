process
    package test is
        signal aaa : bbb;
        signal ccc : ddd := eee;
        signal fff : ggg register;
        signal hhh : iii bus;
        signal jjj : kkk bus := lll;
    end;
begin
end process;
