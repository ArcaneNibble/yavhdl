architecture test of test2 is
    variable foo, foo2 : bar := baz;
begin end;
