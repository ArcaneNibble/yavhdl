entity test is
    type t is range 0 to 16#f.f#e+2;
end;
