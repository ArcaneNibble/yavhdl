entity \test�\ is end;
