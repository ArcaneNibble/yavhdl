entity t__est is end;
